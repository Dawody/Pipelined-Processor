LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.PKG.ALL;

ENTITY MEMORY_BUFFER IS
	PORT (

		D_ALUO1		: IN STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0):=X"0000";
		D_ALUO2		: IN STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0):=X"0000";
		D_MEM		: IN STD_LOGIC_VECTOR(1 DOWNTO 0):="00";		--MEMORY(READ/WRITE)
		D_R_SRC_ADRS	: IN STD_LOGIC_VECTOR(ADDRESS_SIZE-1 DOWNTO 0):="000";
		D_R_DST_ADRS	: IN STD_LOGIC_VECTOR(ADDRESS_SIZE-1 DOWNTO 0):="000";
		D_OPERATION	: IN STD_LOGIC_VECTOR(OPCODE_SIZE-1 DOWNTO 0):="00000";
		D_FLAGS		: IN STD_LOGIC_VECTOR(FLAG_SIZE-1 DOWNTO 0):=X"0";
		D_FE		: IN STD_LOGIC_VECTOR(FLAG_SIZE-1 DOWNTO 0):=X"0";	--FLAGS ENABLE(V-C-N-Z)
		D_A		: IN STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0):=X"0000";
		D_B		: IN STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0):=X"0000";
		
		CLK,RST,ENB	: IN STD_LOGIC;


		Q_ALUO1		:OUT STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0):=X"0000";
		Q_ALUO2		:OUT STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0):=X"0000";
		Q_MEM		:OUT STD_LOGIC_VECTOR(1 DOWNTO 0):="00";		--MEMORY(READ/WRITE)
		Q_R_SRC_ADRS	:OUT STD_LOGIC_VECTOR(ADDRESS_SIZE-1 DOWNTO 0):="000";
		Q_R_DST_ADRS	:OUT STD_LOGIC_VECTOR(ADDRESS_SIZE-1 DOWNTO 0):="000";
		Q_OPERATION	:OUT STD_LOGIC_VECTOR(OPCODE_SIZE-1 DOWNTO 0):="00000";		
		Q_FLAGS		:OUT STD_LOGIC_VECTOR(FLAG_SIZE-1 DOWNTO 0):=X"0";
		Q_FE		:OUT STD_LOGIC_VECTOR(FLAG_SIZE-1 DOWNTO 0):=X"0";	--FLAGS ENABLE(V-C-N-Z)
		Q_A		:OUT STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0):=X"0000";
		Q_B		:OUT STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0):=X"0000"


	);

END ENTITY MEMORY_BUFFER;



ARCHITECTURE MEMORY_BUFFER_ARCH OF MEMORY_BUFFER IS

BEGIN
	PROCESS(CLK,RST,ENB)
		BEGIN
			--IT WILL RESET WHEN I RISE THE RST SIGNAL , IT WILL NOT WAIT TILL THE RISING EDGE.
			--IT WILL RESET ALTHOUGH ENABLE SIGNAL WAS OFF (RST IS POWERFUL THAN EBL)
			IF ((RISING_EDGE(CLK) AND ENB='1') and (RST='1')) THEN
				Q_ALUO1		<= (OTHERS=>'0');
				Q_ALUO2		<= (OTHERS=>'0');
				Q_MEM		<= (OTHERS=>'0');	--MEMORY(READ/WRITE)
				Q_R_SRC_ADRS	<= (OTHERS=>'0');
				Q_R_DST_ADRS	<= (OTHERS=>'0');
				Q_OPERATION	<= (OTHERS=>'0');	
				Q_FLAGS		<= (OTHERS=>'0');
				Q_FE		<= (OTHERS=>'0');	--LAGS ENABLE(V-C-N-Z)
				Q_A		<= (OTHERS=>'0');
				Q_B		<= (OTHERS=>'0');

			ELSIF ((RISING_EDGE(CLK) AND ENB='1')OR(RISING_EDGE(ENB))) THEN
				
				Q_ALUO1		<= D_ALUO1;
				Q_ALUO2		<= D_ALUO2;
				Q_MEM		<= D_MEM;	--MEMORY(READ/WRITE)
				Q_R_SRC_ADRS	<= D_R_SRC_ADRS;
				Q_R_DST_ADRS	<= D_R_DST_ADRS;
				Q_OPERATION	<= D_OPERATION;	
				Q_FLAGS		<= D_FLAGS;
				Q_FE		<= D_FE;	--LAGS ENABLE(V-C-N-Z)
				Q_A		<= D_A;
				Q_B		<= D_B;



			END IF;



	END PROCESS;



END MEMORY_BUFFER_ARCH;