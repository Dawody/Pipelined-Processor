LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL; 

ENTITY FORWARD IS
PORT( OPALU, OPMEM, OPWB: IN std_logic_vector(5 DOWNTO 0);
RSALU, RDALU, RSMEM, RDMEM, RSWB, RDWB: IN std_logic_vector(2 DOWNTO 0);
flags: OUT std_logic_vector(4 DOWNTO 0));
END FORWARD;

ARCHITECTURE struct2 OF FORWARD IS
BEGIN

END struct2;

ENTITY JUMP IS
PORT( tFLAGS: IN std_logic_vector(3 DOWNTO 0);
OPALU: IN std_logic_vector(4 DOWNTO 0);
flu: OUT std_logic);
END JUMP;

ARCHITECTURE struct3 OF JUMP IS
BEGIN

END struct3;