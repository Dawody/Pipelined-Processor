LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.PKG.ALL;



ENTITY FETCH IS 
	PORT(
		ALUO	: IN STD_LOGIC_VECTOR (CELL_SIZE-1 DOWNTO 0);	-- TO BACKWARD THE PC VALUE FROM THE EXECUTION STAGE
		MEMO	: IN STD_LOGIC_VECTOR (CELL_SIZE-1 DOWNTO 0);	-- TO BACKWARD THE PC VALUE FROM THE MEMORY STAGE
		STALL	: IN STD_LOGIC;					-- ENABLE SIGNAL FOR THE PC REGISTER
		INT	: IN STD_LOGIC;					-- INTERRUPT SIGNAL NEEDS PC+1
		FLU1	: IN STD_LOGIC;					-- FLUSH REQUEST COMMING FROM THE JUMP UNIT
		FLU2	: IN STD_LOGIC;					-- FLUSH REQUEST COMMING FROM THE STACK UNIT
		CLK	: IN STD_LOGIC;					-- CLK NEEDED FOR PC REGISTER
		RST,ENB	: IN STD_LOGIC;					-- ACTUALLY, I DON'T NEED THEM NOW. BUT DON'T REMOVE THEM!
		IR	: OUT STD_LOGIC_VECTOR(CELL_SIZE-1 DOWNTO 0);	-- THE INSTRUCTION FORM THE MEMORY
		PC	: OUT STD_LOGIC_VECTOR(CELL_SIZE-1 DOWNTO 0)	-- THE CURRECT PC


	);


END ENTITY FETCH;


ARCHITECTURE FETCH_ARCH OF FETCH IS

------------------------------COMPONENTS----------------------
COMPONENT GENERAL_REGISTER IS
	PORT (
		D		: IN STD_LOGIC_VECTOR (CELL_SIZE-1 DOWNTO 0);
		CLK,RST,ENB	: IN STD_LOGIC;
		Q 		: OUT STD_LOGIC_VECTOR (CELL_SIZE-1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT IR_RAM IS
	PORT (
		ADDRESS		:IN STD_LOGIC_VECTOR(ADDRESS_SIZE-1 DOWNTO 0);
		DATA_OUT 	: OUT STD_LOGIC_VECTOR(CELL_SIZE-1 DOWNTO 0)		
	);
END COMPONENT;

------------------------------SIGNALS------------------------
SIGNAL PC_IN	:STD_LOGIC_VECTOR(CELL_SIZE-1 DOWNTO 0);
SIGNAL PC_OUT	:STD_LOGIC_VECTOR(CELL_SIZE-1 DOWNTO 0);


BEGIN
	RAM	: IR_RAM PORT MAP (ADDRESS => PC_OUT(ADDRESS_SIZE-1 DOWNTO 0) , DATA_OUT => IR);
	REG_PC	: GENERAL_REGISTER PORT MAP (D => PC_IN , CLK => CLK , RST => '0' , ENB => STALL , Q => PC_OUT); --WE CAN IMPROVE THE RESEET SIGNAL TO SUPPORT THE RESET SIGNAL OF THE PROCESSOR (PC <- M[0])


	PC_IN <= ALUO		WHEN FLU1='1'
	ELSE	 MEMO		WHEN FLU2='1' 
	ELSE	 PC_OUT+1;	--ADD THE CASE OF INTERRUPT AND RESET (THEY AFFECT THE PC!)
				--MAKE SURE THAT FLU1 & FLU2 CAN NOT HAPPEN AT THE SAME TIME NEVER!
				--COMP CIRCUIT DO ANY ADDITIONAL FUNCTIONALITY ???



END FETCH_ARCH;