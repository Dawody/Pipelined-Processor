LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.PKG.ALL;



ENTITY FETCH IS 
	PORT(
		ALUO	: IN STD_LOGIC_VECTOR (DATA_SIZE-1 DOWNTO 0);	-- TO BACKWARD THE PC VALUE FROM THE EXECUTION STAGE
		MEMO	: IN STD_LOGIC_VECTOR (DATA_SIZE-1 DOWNTO 0);	-- TO BACKWARD THE PC VALUE FROM THE MEMORY STAGE
		M_1	: IN STD_LOGIC_VECTOR (DATA_SIZE-1 DOWNTO 0);	-- MEM[1] VALUE COMMING FROM THE MEMORY AND NEEDED FOR INTERRUPT CASE (NOTE THAT YOU CAN DO THE SAME IN RESET CASE TO AVOID FLUSHING TWO INSTRUCCTIONS AND WASTING TWO CLK CUCLES!**)		
		STALL	: IN STD_LOGIC;					-- ENABLE SIGNAL FOR THE PC REGISTER
		INT	: IN STD_LOGIC;					-- INTERRUPT SIGNAL NEEDS PC+1
		RESET	: IN STD_LOGIC;					-- RESET THE PROCESSOR!
		FLU1	: IN STD_LOGIC;					-- FLUSH REQUEST COMMING FROM THE JUMP UNIT
		FLU2	: IN STD_LOGIC;					-- FLUSH REQUEST COMMING FROM THE STACK UNIT
		CLK	: IN STD_LOGIC;					-- CLK NEEDED FOR PC REGISTER
		SKIP_IR	: IN STD_LOGIC;					--THIS SIGNAL TO FETCH NEXT IR AS IMMEDIATE OR EFFECTIVE ADDRESS AND SKIP THE CORRESPONDING PC AND FETCH THE CORRECT IR BY INCREMENTING THE PC BY 2
	
		IR	: OUT STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0);	-- THE INSTRUCTION FORM THE MEMORY
		IR_NEXT	: OUT STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0);	--THE NEXT INSTRUCTION THAT MAY BE EFFECTIVE ADDRESS OR IMMEDIATE VALUE NEEDED FOR (LDM,LDD,STD) OPERATIONS	
		PC	: OUT STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0)	-- THE CURRECT PC

	);


END ENTITY FETCH;


ARCHITECTURE FETCH_ARCH OF FETCH IS

------------------------------COMPONENTS----------------------
COMPONENT PC_REGISTER IS
	PORT (
		D		: IN STD_LOGIC_VECTOR (DATA_SIZE-1 DOWNTO 0);
		CLK,RST,ENB	: IN STD_LOGIC;
		FLU		: IN STD_LOGIC;	--THIS SIGNAL RISE ACCORDING TO THE FLUSHES SIGNALS BUT THE ACTUAL PURPOSE FROM THIS SIGNAL IS TO MAKE THE PC REGISTER GET THE NEXT VALUE WITHOUT CLK SIGNAL FOR THIS CLK CYCLE ONLY
		Q 		: OUT STD_LOGIC_VECTOR (DATA_SIZE-1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT IR_RAM IS
	PORT (
		ADDRESS		:IN STD_LOGIC_VECTOR(MEMORY_SIZE-1 DOWNTO 0);
		DATA_OUT 	:OUT STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0);
		NEXT_DATA_OUT	:OUT STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0)		
	);
END COMPONENT;

------------------------------SIGNALS------------------------
SIGNAL PC_IN		:STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0);
SIGNAL PC_OUT		:STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0);
SIGNAL INSTR		:STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0);
SIGNAL NEXT_INSTR	:STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0);
SIGNAL PC_ENB		:STD_LOGIC;
SIGNAL SKIP		:STD_LOGIC;



--------------------------------------------------------------------------------------
BEGIN

	
	RAM	: IR_RAM 	PORT MAP (ADDRESS => PC_OUT(MEMORY_SIZE-1 DOWNTO 0) , DATA_OUT => INSTR , NEXT_DATA_OUT => NEXT_INSTR);
	REG_PC	: PC_REGISTER	PORT MAP (D => PC_IN , CLK => CLK , FLU => SKIP , RST => '0' , ENB => PC_ENB , Q => PC_OUT); --WE CAN IMPROVE THE RESEET SIGNAL TO SUPPORT THE RESET SIGNAL OF THE PROCESSOR (PC <- M[0])

	PC_ENB	<= NOT STALL;
	SKIP 	<= FLU1 OR FLU2 OR SKIP_IR;

	PC_IN <= ALUO		WHEN FLU1='1'	 --LOAD NEW PC VALUE FROM EXECUTION STAGE
	ELSE	 MEMO		WHEN FLU2='1'    --LOAD NEW PC VALUE FROM MEMORY STAGE
	ELSE	 M_1		WHEN INT ='1'    --LOAD NEW PC VALUE FROM M[1] SIGNAL WHEN INTERRUPT
	--ELSE	 PC_OUT+2	WHEN SKIP_IR='1' --THE DECODE STAGE FINDS THAT NEXT IR IS IMMEDIATE OR EFFECTIVE ADRESS SO I NEED TO FETCH THE AFTER NEXT INSTRUCTION AS NEXT IR.
	ELSE	 PC_OUT+1;			 --ORIGINAL CASE

				--MAKE SURE THAT FLU1 & FLU2 CAN NOT HAPPEN AT THE SAME TIME NEVER!**
				--COMP CIRCUIT DO ANY ADDITIONAL FUNCTIONALITY ???**


--------------------------FETCH STAGE OUTPUT-------------------------

	IR 	<= B"11111_110_000_0000_0"	WHEN INT='1'
	ELSE	   B"11110_000_000_0000_0"	WHEN RESET='1'
	ELSE	   INSTR;
	

	IR_NEXT <= NEXT_INSTR;


	PC 	<= PC_OUT		WHEN INT='1' --IN INTERRUPT CASE ONLY I NEED TO SAVE THE CURRENT PC VALUE IN THE REGISTER ; IN OTHER CASES I NEED TO SAVE THE NEXT PC VALUE THAT STAND ON THE ENTRY ON THE REGISTER.
	ELSE	   PC_IN;

	

END FETCH_ARCH;