LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.PKG.ALL;

ENTITY EXECUTE_BUFFER IS
	PORT (

		D_OPERATION	: IN STD_LOGIC_VECTOR(OPCODE_SIZE-1 DOWNTO 0):="00000";
		D_R_SRC_DATA	: IN STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0):=X"0000";
		D_R_DST_DATA	: IN STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0):=X"0000";
		D_FLAGS_DATA	: IN STD_LOGIC_VECTOR(FLAG_SIZE-1 DOWNTO 0):=X"0";
		D_R_SRC_ADRS	: IN STD_LOGIC_VECTOR(ADDRESS_SIZE-1 DOWNTO 0):="000";
		D_R_DST_ADRS	: IN STD_LOGIC_VECTOR(ADDRESS_SIZE-1 DOWNTO 0):="000";
		D_IMMD		: IN STD_LOGIC_VECTOR(3 DOWNTO 0):=X"0";		--IMMEDIATE 4BIT WORKS WITH SHIFT OPERATIONS ONLY
		D_PC		: IN STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0);
		D_MEM_R_W	: IN STD_LOGIC_VECTOR(1 DOWNTO 0):="00";		--MEMORY(READ/WRITE)
		D_FE		: IN STD_LOGIC_VECTOR(FLAG_SIZE-1 DOWNTO 0):=X"0";	--FLAGS ENABLE(V-C-N-Z)
		
		
		CLK,RST,ENB	: IN STD_LOGIC;


		Q_OPERATION	:OUT STD_LOGIC_VECTOR(OPCODE_SIZE-1 DOWNTO 0):="00000";
		Q_R_SRC_DATA	:OUT STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0):=X"0000";
		Q_R_DST_DATA	:OUT STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0):=X"0000";
		Q_FLAGS_DATA	:OUT STD_LOGIC_VECTOR(FLAG_SIZE-1 DOWNTO 0):=X"0";
		Q_R_SRC_ADRS	:OUT STD_LOGIC_VECTOR(ADDRESS_SIZE-1 DOWNTO 0):="000";
		Q_R_DST_ADRS	:OUT STD_LOGIC_VECTOR(ADDRESS_SIZE-1 DOWNTO 0):="000";
		Q_IMMD		:OUT STD_LOGIC_VECTOR(3 DOWNTO 0):=X"0";		--IMMEDIATE 4BIT WORKS WITH SHIFT OPERATIONS ONLY
		Q_PC		:OUT STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0);
		Q_MEM_R_W	:OUT STD_LOGIC_VECTOR(1 DOWNTO 0):="00";		--MEMORY(READ/WRITE)
		Q_FE		:OUT STD_LOGIC_VECTOR(FLAG_SIZE-1 DOWNTO 0):=X"0"	--FLAGS ENABLE(V-C-N-Z)


	);

END ENTITY EXECUTE_BUFFER;



ARCHITECTURE EXECUTE_BUFFER_ARCH OF EXECUTE_BUFFER IS

BEGIN
	PROCESS(CLK,RST,ENB)
		BEGIN
			--IT WILL RESET WHEN I RISE THE RST SIGNAL , IT WILL NOT WAIT TILL THE RISING EDGE.
			--IT WILL RESET ALTHOUGH ENABLE SIGNAL WAS OFF (RST IS POWERFUL THAN EBL)
			IF (RST='1') THEN
				Q_OPERATION	<= (OTHERS=>'0');
				Q_R_SRC_DATA	<= (OTHERS=>'0');
				Q_R_DST_DATA	<= (OTHERS=>'0');
				Q_FLAGS_DATA	<= (OTHERS=>'0');
				Q_R_SRC_ADRS	<= (OTHERS=>'0');
				Q_R_DST_ADRS	<= (OTHERS=>'0');
				Q_IMMD		<= (OTHERS=>'0');
				Q_PC		<= (OTHERS=>'0');
				Q_MEM_R_W	<= (OTHERS=>'0');
				Q_FE		<= (OTHERS=>'0');





			ELSIF ((RISING_EDGE(CLK) AND ENB='1')OR(RISING_EDGE(ENB))) THEN
				Q_OPERATION	<= D_OPERATION;
				Q_R_SRC_DATA	<= D_R_SRC_DATA;
				Q_R_DST_DATA	<= D_R_DST_DATA;
				Q_FLAGS_DATA	<= D_FLAGS_DATA;
				Q_R_SRC_ADRS	<= D_R_SRC_ADRS;
				Q_R_DST_ADRS	<= D_R_DST_ADRS;
				Q_IMMD		<= D_IMMD;
				Q_PC		<= D_PC;
				Q_MEM_R_W	<= D_MEM_R_W;
				Q_FE		<= D_FE;

			END IF;



	END PROCESS;



END EXECUTE_BUFFER_ARCH;