LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.PKG.ALL;




ENTITY IR_RAM IS
	--GENERIC (ADDRESS_SIZE : INTEGER :=11; CELL_SIZE : INTEGER := 16*2);	--11BIT FOR MEMORY ADDRESS_SIZE PROVIDES 2K BIT MEMORY --16*2 : I ALLWAYS READ & WRITE 2 CELLS BUT I MAYBE WANT TO READ 1 CELL IN THIS CASE MDR WILL HANDLE IT
	PORT (
		ADDRESS		:IN STD_LOGIC_VECTOR(MEMORY_SIZE-1 DOWNTO 0);
		DATA_OUT 	:OUT STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0);
		NEXT_DATA_OUT	:OUT STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0)		
	);
END ENTITY IR_RAM;
		

ARCHITECTURE IR_RAM_ARCH OF IR_RAM IS

	TYPE RAM_TYPE IS ARRAY(0 TO 1024) OF std_logic_vector(DATA_SIZE-1 DOWNTO 0);
	SIGNAL MEMORY : RAM_TYPE ;
	
	BEGIN
		DATA_OUT 	<= MEMORY(to_integer(unsigned(ADDRESS)));
		NEXT_DATA_OUT	<= MEMORY(TO_INTEGER(UNSIGNED(ADDRESS+1)));
		

END IR_RAM_ARCH;
