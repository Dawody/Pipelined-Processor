LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.PKG.ALL;



ENTITY FETCH IS 
	PORT(
		ALUO	: IN STD_LOGIC_VECTOR (DATA_SIZE-1 DOWNTO 0);	-- TO BACKWARD THE PC VALUE FROM THE EXECUTION STAGE
		MEMO	: IN STD_LOGIC_VECTOR (DATA_SIZE-1 DOWNTO 0);	-- TO BACKWARD THE PC VALUE FROM THE MEMORY STAGE
		M_1	: IN STD_LOGIC_VECTOR (DATA_SIZE-1 DOWNTO 0);	-- MEM[1] VALUE COMMING FROM THE MEMORY AND NEEDED FOR INTERRUPT CASE (NOTE THAT YOU CAN DO THE SAME IN RESET CASE TO AVOID FLUSHING TWO INSTRUCCTIONS AND WASTING TWO CLK CUCLES!**)		
		STALL	: IN STD_LOGIC;					-- ENABLE SIGNAL FOR THE PC REGISTER
		INT	: IN STD_LOGIC;					-- INTERRUPT SIGNAL NEEDS PC+1
		FLU1	: IN STD_LOGIC;					-- FLUSH REQUEST COMMING FROM THE JUMP UNIT
		FLU2	: IN STD_LOGIC;					-- FLUSH REQUEST COMMING FROM THE STACK UNIT
		CLK	: IN STD_LOGIC;					-- CLK NEEDED FOR PC REGISTER
		RST,ENB	: IN STD_LOGIC;					-- ACTUALLY, I DON'T NEED THEM NOW. BUT DON'T REMOVE THEM!
		IR	: OUT STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0);	-- THE INSTRUCTION FORM THE MEMORY
		PC	: OUT STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0)	-- THE CURRECT PC

	);


END ENTITY FETCH;


ARCHITECTURE FETCH_ARCH OF FETCH IS

------------------------------COMPONENTS----------------------
COMPONENT PC_REGISTER IS
	PORT (
		D		: IN STD_LOGIC_VECTOR (DATA_SIZE-1 DOWNTO 0);
		CLK,RST,ENB	: IN STD_LOGIC;
		Q 		: OUT STD_LOGIC_VECTOR (DATA_SIZE-1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT IR_RAM IS
	PORT (
		ADDRESS		:IN STD_LOGIC_VECTOR(MEMORY_SIZE-1 DOWNTO 0);
		DATA_OUT 	: OUT STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0)		
	);
END COMPONENT;

------------------------------SIGNALS------------------------
SIGNAL PC_IN	:STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0);
SIGNAL PC_OUT	:STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0);
SIGNAL INSTR	:STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0);
SIGNAL PC_ENB	:STD_LOGIC;


--------------------------------------------------------------------------------------
BEGIN

	
	RAM	: IR_RAM 	PORT MAP (ADDRESS => PC_OUT(MEMORY_SIZE-1 DOWNTO 0) , DATA_OUT => INSTR);
	REG_PC	: PC_REGISTER	PORT MAP (D => PC_IN , CLK => CLK , RST => '0' , ENB => PC_ENB , Q => PC_OUT); --WE CAN IMPROVE THE RESEET SIGNAL TO SUPPORT THE RESET SIGNAL OF THE PROCESSOR (PC <- M[0])

	PC_ENB <= NOT STALL;

	PC_IN <= ALUO		WHEN FLU1='1' --LOAD NEW PC VALUE FROM EXECUTION STAGE
	ELSE	 MEMO		WHEN FLU2='1' --LOAD NEW PC VALUE FROM MEMORY STAGE
	ELSE	 M_1		WHEN INT ='1' --LOAD NEW PC VALUE FROM M[1] SIGNAL WHEN INTERRUPT
	ELSE	 PC_OUT+1;	
				--MAKE SURE THAT FLU1 & FLU2 CAN NOT HAPPEN AT THE SAME TIME NEVER!**
				--COMP CIRCUIT DO ANY ADDITIONAL FUNCTIONALITY ???**


--------------------------FETCH STAGE OUTPUT-------------------------

	IR <=	INSTR		WHEN INT='0'
	ELSE	"1111111111111111";	--RESET??**
					

	PC <=	PC_OUT		WHEN INT='1' --IN INTERRUPT CASE ONLY I NEED TO SAVE THE CURRENT PC VALUE IN THE REGISTER ; IN OTHER CASES I NEED TO SAVE THE NEXT PC VALUE THAT STAND ON THE ENTRY ON THE REGISTER.
	ELSE	PC_IN;

	

END FETCH_ARCH;